magic
tech sky130A
magscale 1 2
timestamp 1729046266
<< error_p >>
rect 79 515 239 549
rect 298 515 335 532
rect 299 514 335 515
rect 299 478 371 514
rect 316 453 389 478
rect -17 79 19 453
rect 129 447 189 453
rect 129 413 177 447
rect 299 444 389 453
rect 448 444 608 478
rect 129 407 189 413
rect 97 178 133 354
rect 143 178 144 365
rect 174 354 175 365
rect 185 178 221 354
rect 141 85 177 119
rect 299 79 388 444
rect 498 376 558 382
rect 498 342 546 376
rect 498 336 558 342
rect 466 116 502 292
rect 512 116 513 303
rect 543 292 544 303
rect 554 116 590 292
rect 79 -17 239 17
rect 316 -17 388 79
rect 498 66 558 72
rect 498 32 546 66
rect 498 26 558 32
rect 668 26 704 382
rect 316 -53 371 -17
rect 448 -70 608 -36
use oscillator  x1
timestamp 1729046265
transform 1 0 53 0 1 2106
box -106 -2212 687 200
<< end >>
