magic
tech sky130A
magscale 1 2
timestamp 1729443144
<< error_p >>
rect 98 1809 123 1843
rect 132 1785 157 1809
rect 331 1798 556 1809
rect 342 1786 556 1798
rect 331 1785 556 1786
rect 132 1775 556 1785
rect 600 1778 800 1790
rect 55 441 70 1775
rect 89 494 123 1775
rect 178 1723 242 1741
rect 296 1731 330 1741
rect 522 1735 556 1775
rect 575 1753 834 1756
rect 847 1753 899 1756
rect 522 1731 542 1735
rect 296 1723 343 1731
rect 178 1707 254 1723
rect 284 1707 343 1723
rect 380 1707 427 1731
rect 196 1673 427 1707
rect 150 1626 157 1630
rect 174 1626 184 1630
rect 196 1626 254 1673
rect 284 1626 342 1673
rect 138 1331 190 1626
rect 202 1356 242 1626
rect 202 1343 248 1356
rect 202 1331 218 1343
rect 226 1331 248 1343
rect 254 1331 276 1356
rect 296 1343 330 1626
rect 397 1614 442 1625
rect 408 1331 442 1614
rect 522 1331 556 1731
rect 575 1722 968 1753
rect 1018 1722 1033 1790
rect 1060 1722 1095 1756
rect 138 1284 289 1331
rect 396 1284 454 1331
rect 138 1226 190 1284
rect 192 1250 289 1284
rect 358 1250 454 1284
rect 192 1244 218 1250
rect 192 1235 196 1244
rect 396 1234 454 1250
rect 439 1226 454 1234
rect 522 1327 542 1331
rect 522 1234 556 1327
rect 150 1222 157 1226
rect 158 1222 184 1226
rect 522 1223 533 1234
rect 300 1129 396 1170
rect 522 1128 533 1139
rect 541 1128 556 1234
rect 371 1112 420 1118
rect 342 1111 430 1112
rect 383 1105 418 1111
rect 284 1080 430 1105
rect 342 1078 430 1080
rect 364 1077 371 1078
rect 284 1071 371 1077
rect 254 1069 396 1071
rect 196 1044 396 1069
rect 196 1037 380 1044
rect 522 1035 556 1128
rect 208 1031 242 1035
rect 296 1031 330 1035
rect 522 1031 542 1035
rect 150 990 157 994
rect 174 990 184 994
rect 196 990 254 1031
rect 284 990 342 1031
rect 138 631 190 990
rect 202 643 242 990
rect 296 643 330 990
rect 397 978 442 989
rect 202 631 218 643
rect 408 631 442 978
rect 522 631 556 1031
rect 138 590 289 631
rect 311 590 454 631
rect 522 627 542 631
rect 146 584 218 590
rect 408 586 442 590
rect 146 577 242 584
rect 358 580 480 584
rect 374 577 480 580
rect 146 550 258 577
rect 342 564 480 577
rect 342 552 476 564
rect 342 550 430 552
rect 146 549 196 550
rect 364 549 371 550
rect 196 528 292 543
rect 308 528 396 543
rect 196 509 396 528
rect 522 534 556 627
rect 522 528 533 534
rect 541 528 556 534
rect 522 503 556 528
rect 541 494 556 503
rect 575 494 609 1722
rect 793 1671 806 1688
rect 812 1670 859 1701
rect 900 1688 946 1701
rect 900 1670 953 1688
rect 800 1660 859 1670
rect 765 1654 859 1660
rect 888 1654 953 1670
rect 751 1620 953 1654
rect 1027 1627 1052 1722
rect 800 1573 858 1620
rect 888 1601 935 1620
rect 888 1573 940 1601
rect 947 1573 968 1577
rect 678 1561 723 1572
rect 689 1331 723 1561
rect 812 1343 846 1573
rect 900 1343 940 1573
rect 677 1284 736 1331
rect 784 1284 831 1331
rect 913 1330 940 1343
rect 941 1561 968 1573
rect 941 1330 972 1561
rect 677 1250 831 1284
rect 853 1283 981 1330
rect 677 1173 735 1250
rect 900 1249 981 1283
rect 935 1234 972 1249
rect 947 1211 972 1234
rect 1018 1173 1052 1627
rect 725 1112 919 1126
rect 616 1092 919 1112
rect 616 1078 784 1092
rect 816 1076 930 1092
rect 812 1031 846 1052
rect 900 1031 953 1052
rect 800 1018 859 1031
rect 888 1018 953 1031
rect 751 984 953 1018
rect 1027 991 1052 1173
rect 800 937 858 984
rect 888 937 935 984
rect 678 925 723 936
rect 689 631 723 925
rect 812 643 846 937
rect 900 643 934 937
rect 913 634 934 643
rect 947 925 968 941
rect 947 634 972 925
rect 913 631 940 634
rect 941 631 972 634
rect 677 584 736 631
rect 784 584 831 631
rect 853 584 981 631
rect 677 550 831 584
rect 900 550 981 584
rect 677 537 735 550
rect 935 549 972 550
rect 935 548 965 549
rect 935 537 993 548
rect 1018 537 1052 991
rect 717 494 953 524
rect 89 490 992 494
rect 89 460 957 490
rect 1027 460 1052 537
rect 55 426 522 441
rect 541 407 556 460
rect 575 407 609 460
rect 1061 426 1095 1722
rect 575 373 590 407
rect 1080 354 1095 426
rect 1114 1669 1149 1703
rect 1599 1669 1634 1703
rect 1114 354 1148 1669
rect 1600 1650 1634 1669
rect 1114 320 1129 354
rect 1619 301 1634 1650
rect 1653 1616 1688 1650
rect 1968 1616 2003 1650
rect 1653 301 1687 1616
rect 1969 1597 2003 1616
rect 1799 1548 1857 1554
rect 1799 1514 1811 1548
rect 1799 1508 1857 1514
rect 1799 1020 1857 1026
rect 1799 986 1811 1020
rect 1799 980 1857 986
rect 1799 912 1857 918
rect 1799 878 1811 912
rect 1799 872 1857 878
rect 1799 384 1857 390
rect 1799 350 1811 384
rect 1799 344 1857 350
rect 1653 267 1668 301
rect 1988 248 2003 1597
rect 2022 1563 2057 1597
rect 2022 248 2056 1563
rect 2022 214 2037 248
rect 8831 2077 8841 2156
rect 8773 1973 8784 1984
rect 8796 1973 8807 1984
rect 8773 1878 8784 1889
rect 8796 1878 8807 1889
rect 8733 1828 8752 1862
rect 8733 1500 8752 1534
rect 8831 1577 8841 1785
rect 8773 1473 8784 1484
rect 8796 1473 8807 1484
rect 8773 1379 8784 1390
rect 8796 1379 8807 1390
rect 8733 1329 8752 1363
rect 8733 1082 8759 1121
rect 8733 1001 8752 1035
rect 8831 1197 8841 1286
rect 9131 1197 9165 1981
rect 10019 1929 10054 1963
rect 10020 1910 10054 1929
rect 9850 1861 9908 1867
rect 9850 1827 9862 1861
rect 9850 1821 9908 1827
rect 9850 1533 9908 1539
rect 9850 1499 9862 1533
rect 9850 1493 9908 1499
rect 9850 1425 9908 1431
rect 9850 1391 9862 1425
rect 9850 1385 9908 1391
rect 9077 1163 9165 1197
rect 9211 1163 9246 1197
rect 8964 1129 8977 1133
rect 8952 1097 8977 1129
rect 9031 1111 9077 1142
rect 8952 1082 8986 1097
rect 8989 1082 9002 1095
rect 9077 1094 9099 1095
rect 8826 1069 8841 1082
rect 8939 1073 9015 1082
rect 9019 1073 9069 1082
rect 8939 1069 9069 1073
rect 8807 1001 8819 1035
rect 8773 974 8784 985
rect 8773 880 8784 891
rect 8792 880 8807 985
rect 8733 830 8735 864
rect 8733 502 8752 536
rect 8826 985 8853 1069
rect 8939 1061 9070 1069
rect 8990 1055 9061 1061
rect 8975 1035 9033 1041
rect 9131 1036 9165 1163
rect 9212 1144 9246 1163
rect 8936 1027 9037 1035
rect 8936 1014 8986 1027
rect 8956 1002 8971 1014
rect 8949 985 8971 1002
rect 8987 1023 9021 1027
rect 8987 1014 9012 1023
rect 9131 1014 9166 1036
rect 9021 1001 9068 1014
rect 8826 880 8860 985
rect 8949 963 8980 985
rect 8959 902 8980 963
rect 8949 880 8980 902
rect 8807 830 8819 864
rect 8826 837 8853 880
rect 8949 837 8971 880
rect 8826 783 8860 837
rect 8928 814 8971 837
rect 8987 870 9008 995
rect 9021 830 9068 911
rect 8989 824 9019 830
rect 9098 826 9131 860
rect 8987 814 9019 824
rect 9144 826 9166 1014
rect 8940 810 8974 814
rect 8943 783 8977 787
rect 8987 786 9008 814
rect 9031 783 9065 801
rect 8943 776 8986 783
rect 8952 768 8986 776
rect 8952 699 8977 768
rect 8989 733 9002 767
rect 9077 733 9099 767
rect 9062 706 9077 717
rect 8964 693 8977 699
rect 8952 632 8977 693
rect 9031 675 9077 706
rect 8874 583 8877 632
rect 8931 606 8986 632
rect 8906 583 8986 606
rect 8989 625 9002 659
rect 9077 625 9099 659
rect 8989 583 9019 625
rect 9131 600 9140 632
rect 8807 502 8819 536
rect 8773 464 8807 486
rect 8826 464 8860 583
rect 8940 582 8943 583
rect 9064 579 9065 583
rect 9098 578 9099 582
rect 8934 555 8980 578
rect 9092 566 9099 578
rect 9131 578 9166 600
rect 9092 555 9098 566
rect 8940 464 8974 498
rect 9098 464 9131 498
rect 9144 524 9166 578
rect 8733 430 8928 464
rect 9212 430 9219 1144
rect 8773 344 8807 430
rect 8792 248 8807 344
rect 8826 248 8860 430
rect 8826 214 8841 248
rect 9231 195 9246 1144
rect 9265 1110 9300 1144
rect 9265 195 9299 1110
rect 9265 161 9280 195
rect 9670 142 9685 1144
rect 9704 142 9738 1198
rect 9850 1097 9908 1103
rect 9850 1063 9862 1097
rect 9850 1057 9908 1063
rect 9850 989 9908 995
rect 9850 955 9862 989
rect 9850 949 9908 955
rect 9850 661 9908 667
rect 9850 627 9862 661
rect 9850 621 9908 627
rect 9850 553 9908 559
rect 9850 519 9862 553
rect 9850 513 9908 519
rect 9850 225 9908 231
rect 9850 191 9862 225
rect 9850 185 9908 191
rect 9704 108 9719 142
rect 10039 89 10054 1910
rect 10073 1876 10108 1910
rect 10073 89 10107 1876
rect 10219 1808 10277 1814
rect 10219 1774 10231 1808
rect 10219 1768 10277 1774
rect 10219 1480 10277 1486
rect 10219 1446 10231 1480
rect 10219 1440 10277 1446
rect 10219 1372 10277 1378
rect 10219 1338 10231 1372
rect 10219 1332 10277 1338
rect 10219 1044 10277 1050
rect 10219 1010 10231 1044
rect 10219 1004 10277 1010
rect 10219 936 10277 942
rect 10219 902 10231 936
rect 10219 896 10277 902
rect 10219 608 10277 614
rect 10219 574 10231 608
rect 10219 568 10277 574
rect 10219 500 10277 506
rect 10219 466 10231 500
rect 10219 460 10277 466
rect 10219 172 10277 178
rect 10219 138 10231 172
rect 10219 132 10277 138
rect 10073 55 10088 89
<< error_s >>
rect 7571 2228 7597 2262
rect 7663 2228 7697 2285
rect 7751 2228 7785 2285
rect 7863 2228 7867 2262
rect 7605 2194 7631 2228
rect 7651 2194 7797 2228
rect 7851 2194 7929 2228
rect 6035 1963 6070 1997
rect 6036 1944 6070 1963
rect 6055 1901 6070 1944
rect 2507 1563 2542 1597
rect 2508 1544 2542 1563
rect 2527 195 2542 1544
rect 2561 1510 2596 1544
rect 2876 1510 2911 1544
rect 4206 1527 4241 1561
rect 2561 195 2595 1510
rect 2877 1491 2911 1510
rect 4207 1508 4241 1527
rect 2707 1442 2765 1448
rect 2707 1408 2719 1442
rect 2707 1402 2765 1408
rect 2707 914 2765 920
rect 2707 880 2719 914
rect 2707 874 2765 880
rect 2707 806 2765 812
rect 2707 772 2719 806
rect 2707 766 2765 772
rect 2707 278 2765 284
rect 2707 244 2719 278
rect 2707 238 2765 244
rect 2561 161 2576 195
rect 2896 142 2911 1491
rect 2930 1457 2965 1491
rect 3245 1457 3280 1491
rect 2930 142 2964 1457
rect 3246 1438 3280 1457
rect 3076 1389 3134 1395
rect 3076 1355 3088 1389
rect 3076 1349 3134 1355
rect 3076 861 3134 867
rect 3076 827 3088 861
rect 3076 821 3134 827
rect 3076 753 3134 759
rect 3076 719 3088 753
rect 3076 713 3134 719
rect 3076 225 3134 231
rect 3076 191 3088 225
rect 3076 185 3134 191
rect 2930 108 2945 142
rect 3265 89 3280 1438
rect 3299 1404 3334 1438
rect 3299 89 3333 1404
rect 3721 1398 3755 1465
rect 3897 1459 4065 1492
rect 4226 1465 4241 1508
rect 4207 1458 4241 1465
rect 4260 1474 4746 1508
rect 4260 1458 4294 1474
rect 3870 1455 4962 1458
rect 3870 1447 5053 1455
rect 3881 1441 5053 1447
rect 3769 1424 5053 1441
rect 3769 1398 3772 1424
rect 3445 1336 3503 1342
rect 3445 1302 3457 1336
rect 3445 1296 3503 1302
rect 3445 808 3503 814
rect 3445 774 3457 808
rect 3445 768 3503 774
rect 3445 700 3503 706
rect 3445 666 3457 700
rect 3445 660 3503 666
rect 3721 291 3772 1398
rect 3835 1390 3869 1391
rect 4071 1387 4127 1393
rect 3823 987 3826 1387
rect 3835 1309 3881 1375
rect 3917 1359 3955 1387
rect 4071 1359 4139 1387
rect 3883 1325 3955 1359
rect 4089 1325 4165 1359
rect 4089 1315 4139 1325
rect 3835 1275 3869 1309
rect 4059 1287 4077 1291
rect 4087 1287 4139 1315
rect 4059 1286 4083 1287
rect 3835 999 3873 1275
rect 3839 983 3873 999
rect 3881 987 3884 1286
rect 3916 1275 3961 1286
rect 4032 1275 4083 1286
rect 3927 987 3961 1275
rect 4043 987 4083 1275
rect 4087 999 4127 1287
rect 4087 987 4123 999
rect 3839 899 3879 983
rect 3881 955 3885 987
rect 3881 949 3907 955
rect 3915 949 3973 987
rect 3881 915 3973 949
rect 3881 909 3907 915
rect 3881 899 3885 909
rect 3915 899 3973 915
rect 3847 887 3879 899
rect 3847 883 3873 887
rect 3885 861 3915 899
rect 3958 887 3973 899
rect 4031 983 4083 987
rect 4093 983 4111 987
rect 4031 915 4099 983
rect 4031 899 4081 915
rect 4031 887 4046 899
rect 4055 815 4081 841
rect 3881 807 3996 815
rect 4009 807 4081 815
rect 3885 801 3996 805
rect 4009 801 4077 805
rect 3847 777 3874 781
rect 3928 777 3962 781
rect 4043 777 4077 781
rect 4089 777 4123 899
rect 3847 773 3886 777
rect 3866 769 3886 773
rect 3916 769 3974 777
rect 4031 769 4089 777
rect 4093 769 4111 773
rect 3823 369 3826 769
rect 3866 765 3885 769
rect 3917 765 3962 769
rect 4032 768 4123 769
rect 4032 765 4127 768
rect 3840 762 3885 765
rect 3840 757 3874 762
rect 3835 389 3874 757
rect 3881 389 3885 762
rect 3928 389 3962 765
rect 4043 389 4077 765
rect 4081 762 4127 765
rect 4089 389 4127 762
rect 3835 381 3869 389
rect 4059 384 4083 389
rect 4087 384 4127 389
rect 4059 381 4127 384
rect 4059 377 4123 381
rect 3846 373 3956 377
rect 4059 373 4077 377
rect 3835 369 3956 373
rect 4081 369 4139 377
rect 3835 365 3869 369
rect 4089 365 4127 369
rect 4089 345 4123 365
rect 3874 341 3903 345
rect 4089 341 4161 345
rect 4089 339 4123 341
rect 3868 331 3931 339
rect 4089 331 4161 339
rect 3884 305 4081 331
rect 3897 297 4081 305
rect 3738 278 3772 291
rect 4089 289 4123 331
rect 4207 289 4241 1424
rect 4207 278 4218 289
rect 4226 252 4241 289
rect 4260 252 4294 1424
rect 4765 1412 4780 1424
rect 4420 1390 4620 1406
rect 4439 1372 4620 1390
rect 4474 1366 4616 1372
rect 4370 1334 4420 1364
rect 4502 1359 4644 1365
rect 4473 1338 4654 1359
rect 4514 1334 4632 1338
rect 4644 1334 4654 1338
rect 4362 1314 4420 1334
rect 4489 1325 4678 1334
rect 4620 1319 4678 1325
rect 4301 883 4328 1291
rect 4340 906 4341 1287
rect 4362 1275 4414 1314
rect 4427 1287 4442 1291
rect 4620 1287 4673 1319
rect 4685 1287 4700 1291
rect 4421 1286 4442 1287
rect 4420 1275 4461 1286
rect 4362 934 4408 1275
rect 4427 934 4461 1275
rect 4632 1043 4672 1287
rect 4679 1275 4700 1287
rect 4679 1043 4704 1275
rect 4632 952 4666 1043
rect 4685 952 4704 1043
rect 4632 946 4672 952
rect 4651 934 4672 946
rect 4393 930 4408 934
rect 4415 896 4473 934
rect 4604 896 4642 934
rect 4651 930 4666 934
rect 4679 908 4704 952
rect 4679 906 4700 908
rect 4685 899 4700 906
rect 4415 887 4642 896
rect 4436 883 4604 887
rect 4712 883 4719 1291
rect 4721 887 4731 1287
rect 4436 877 4620 883
rect 4424 862 4620 877
rect 4424 856 4616 862
rect 4502 849 4644 855
rect 4396 828 4461 849
rect 4473 828 4654 849
rect 4514 822 4632 828
rect 4396 815 4426 822
rect 4473 815 4654 822
rect 4502 809 4644 815
rect 4436 794 4495 799
rect 4424 787 4426 794
rect 4436 788 4616 794
rect 4301 770 4328 781
rect 4427 777 4436 788
rect 4439 781 4620 788
rect 4476 777 4604 781
rect 4301 744 4347 770
rect 4415 762 4642 777
rect 4420 754 4642 762
rect 4301 716 4353 744
rect 4393 716 4408 720
rect 4420 716 4473 754
rect 4685 744 4700 754
rect 4679 742 4700 744
rect 4651 716 4666 720
rect 4301 373 4328 716
rect 4340 389 4353 716
rect 4340 377 4341 389
rect 4362 377 4414 716
rect 4421 389 4461 716
rect 4651 715 4672 716
rect 4621 704 4672 715
rect 4421 377 4442 389
rect 4632 377 4672 704
rect 4679 389 4704 742
rect 4679 377 4700 389
rect 4368 365 4381 377
rect 4362 361 4381 365
rect 4362 350 4377 361
rect 4389 351 4414 377
rect 4393 350 4414 351
rect 4362 316 4420 350
rect 4370 300 4420 316
rect 4427 288 4442 377
rect 4620 373 4673 377
rect 4685 373 4700 377
rect 4712 373 4719 781
rect 4721 377 4731 777
rect 4620 362 4691 373
rect 4598 339 4691 362
rect 4489 328 4691 339
rect 4489 316 4678 328
rect 4514 312 4632 316
rect 4473 305 4654 312
rect 4502 299 4644 305
rect 4436 284 4604 286
rect 4436 278 4616 284
rect 4432 252 4436 278
rect 4439 271 4620 278
rect 4476 267 4604 271
rect 4746 252 4780 1412
rect 4799 1421 4834 1424
rect 4895 1421 5053 1424
rect 5114 1421 5149 1455
rect 4799 1287 4833 1421
rect 5115 1402 5149 1421
rect 4988 1387 5022 1400
rect 4917 1291 4922 1365
rect 4988 1359 5025 1387
rect 4945 1353 5025 1359
rect 4945 1325 4957 1353
rect 4941 1319 4957 1325
rect 4988 1319 5025 1353
rect 4945 1313 5007 1319
rect 4988 1303 5007 1313
rect 4788 887 4834 1287
rect 4907 1285 4922 1291
rect 4888 1269 4922 1275
rect 4967 1269 5022 1303
rect 4888 899 4947 1269
rect 4913 893 4947 899
rect 4988 893 5056 1269
rect 4799 777 4833 887
rect 4988 877 5022 893
rect 4988 849 5025 877
rect 4945 843 5025 849
rect 4945 809 4957 843
rect 4988 809 5025 843
rect 4945 803 5007 809
rect 4988 793 5007 803
rect 4988 782 4999 793
rect 4787 377 4834 777
rect 4988 769 5022 782
rect 4887 670 4933 765
rect 4988 741 5025 769
rect 4945 735 5025 741
rect 4941 701 4971 735
rect 4988 701 5025 735
rect 4945 695 5007 701
rect 4988 685 5007 695
rect 4887 667 4927 670
rect 4887 651 4921 667
rect 4967 651 5022 685
rect 4887 389 4947 651
rect 4913 377 4947 389
rect 4799 252 4833 377
rect 4875 305 4877 339
rect 4879 305 4893 339
rect 4901 306 4947 377
rect 4901 263 4959 306
rect 4988 278 5056 651
rect 4913 259 4947 263
rect 4923 252 4962 259
rect 4988 252 5022 278
rect 3798 218 5022 252
rect 3817 195 4145 218
rect 4226 195 4241 218
rect 4260 195 4294 218
rect 3445 172 3503 178
rect 3445 138 3457 172
rect 4260 161 4275 195
rect 4765 142 4780 218
rect 4799 142 4833 218
rect 4945 191 4957 218
rect 4945 185 5003 191
rect 3445 132 3503 138
rect 4799 108 4814 142
rect 5134 89 5149 1402
rect 5168 1368 5203 1402
rect 5590 1386 5624 1901
rect 5766 1477 5894 1480
rect 6036 1447 6070 1901
rect 6089 1910 6124 1944
rect 6036 1446 6087 1447
rect 6089 1446 6123 1910
rect 6231 1446 6427 1458
rect 6535 1446 6569 1848
rect 6957 1446 6991 1742
rect 7059 1464 7103 1500
rect 7071 1460 7083 1464
rect 5638 1412 6992 1446
rect 7037 1426 7049 1446
rect 5638 1405 5641 1412
rect 5704 1405 5738 1409
rect 5922 1405 5956 1409
rect 5692 1403 5750 1405
rect 5692 1399 5779 1403
rect 5673 1387 5779 1399
rect 5910 1387 5968 1405
rect 5168 89 5202 1368
rect 5314 1300 5372 1306
rect 5314 1266 5326 1300
rect 5314 1260 5372 1266
rect 5314 790 5372 796
rect 5314 756 5326 790
rect 5314 750 5372 756
rect 5314 682 5372 688
rect 5314 648 5326 682
rect 5314 642 5372 648
rect 5590 291 5641 1386
rect 5673 1381 5738 1387
rect 5741 1381 5779 1387
rect 5673 1365 5779 1381
rect 5922 1377 5968 1387
rect 5692 1331 5779 1365
rect 5910 1361 5968 1377
rect 5692 1315 5750 1331
rect 5857 1327 5968 1361
rect 5692 1300 5738 1315
rect 5692 1205 5695 1300
rect 5704 1277 5738 1300
rect 5910 1289 5968 1327
rect 6036 1293 6070 1412
rect 5704 1217 5741 1277
rect 5692 833 5695 987
rect 5707 975 5741 1217
rect 5750 1205 5752 1288
rect 5784 1277 5829 1288
rect 5795 1205 5829 1277
rect 5922 1217 5956 1289
rect 5750 1167 5753 1205
rect 5783 1167 5841 1205
rect 5894 1167 5932 1205
rect 5750 1133 5932 1167
rect 5750 1117 5753 1133
rect 5783 1117 5841 1133
rect 5795 1075 5833 1097
rect 5704 901 5741 975
rect 5750 1059 5753 1075
rect 5783 1059 5841 1075
rect 5894 1059 5932 1097
rect 5750 1025 5932 1059
rect 5750 987 5753 1025
rect 5783 987 5841 1025
rect 5750 901 5752 987
rect 5795 901 5829 987
rect 5911 975 5956 986
rect 5704 833 5738 901
rect 5922 889 5956 975
rect 5910 851 5968 889
rect 5857 833 5968 851
rect 5692 787 5750 833
rect 5753 787 5783 833
rect 5841 787 5968 833
rect 6036 885 6087 1293
rect 6036 817 6070 885
rect 5738 783 5741 787
rect 5716 779 5741 783
rect 5795 779 5829 783
rect 6036 779 6041 817
rect 6055 783 6070 817
rect 6055 779 6087 783
rect 5701 759 5772 779
rect 5692 378 5695 569
rect 5707 557 5741 759
rect 5750 749 5753 759
rect 5783 749 5841 779
rect 5894 749 5932 779
rect 5750 715 5932 749
rect 5750 699 5753 715
rect 5783 699 5841 715
rect 5795 657 5833 679
rect 5704 391 5741 557
rect 5750 641 5753 657
rect 5783 641 5841 657
rect 5894 641 5932 679
rect 5750 607 5932 641
rect 5750 569 5753 607
rect 5783 569 5841 607
rect 5750 391 5752 569
rect 5795 391 5829 569
rect 5911 557 5956 568
rect 5704 381 5738 391
rect 5922 381 5956 557
rect 5692 369 5779 378
rect 5819 369 5968 379
rect 6036 375 6087 779
rect 5704 365 5707 369
rect 5922 365 5956 369
rect 5726 346 5747 365
rect 5695 341 5702 346
rect 5691 331 5707 340
rect 5726 300 5753 346
rect 5888 341 5990 347
rect 5757 337 5784 340
rect 5754 331 5784 337
rect 5857 331 6025 341
rect 5754 307 6025 331
rect 6036 307 6070 375
rect 5754 297 5894 307
rect 5754 291 5781 297
rect 6036 293 6041 307
rect 6055 293 6070 307
rect 6036 291 6070 293
rect 5607 285 5641 291
rect 6036 280 6047 291
rect 6055 260 6070 291
rect 6055 259 6087 260
rect 6089 259 6123 1412
rect 6265 1395 6296 1399
rect 6360 1395 6393 1399
rect 6249 1390 6409 1395
rect 6253 1384 6298 1390
rect 6358 1384 6405 1390
rect 6169 1361 6271 1374
rect 6387 1367 6489 1374
rect 6386 1361 6489 1367
rect 6535 1361 6569 1412
rect 6215 1356 6299 1361
rect 6357 1356 6443 1361
rect 6227 1352 6258 1356
rect 6398 1352 6431 1356
rect 6191 1327 6321 1352
rect 6373 1327 6467 1352
rect 6191 1289 6249 1327
rect 6409 1289 6467 1327
rect 6535 1311 6557 1361
rect 6561 1311 6569 1343
rect 6203 1164 6237 1289
rect 6300 1277 6345 1288
rect 6311 1152 6345 1277
rect 6421 1164 6455 1289
rect 6299 1114 6357 1152
rect 6393 1114 6431 1152
rect 6265 1080 6431 1114
rect 6299 1064 6357 1080
rect 6311 1022 6349 1044
rect 6299 1006 6357 1022
rect 6393 1006 6431 1044
rect 6265 972 6431 1006
rect 6299 934 6357 972
rect 6192 922 6237 933
rect 6203 889 6237 922
rect 6311 901 6345 934
rect 6410 922 6455 933
rect 6421 889 6455 922
rect 6535 889 6569 1311
rect 6923 1055 6949 1331
rect 6588 1021 6949 1055
rect 6191 851 6249 889
rect 6283 851 6321 889
rect 6409 851 6467 889
rect 6191 817 6321 851
rect 6373 817 6467 851
rect 6191 779 6249 817
rect 6409 779 6467 817
rect 6535 885 6557 889
rect 6203 746 6237 779
rect 6300 767 6345 778
rect 6311 734 6345 767
rect 6421 746 6455 779
rect 6299 696 6357 734
rect 6393 696 6431 734
rect 6265 662 6431 696
rect 6299 646 6357 662
rect 6311 604 6349 626
rect 6299 588 6357 604
rect 6393 588 6431 626
rect 6265 554 6431 588
rect 6299 516 6357 554
rect 6192 504 6237 515
rect 6203 379 6237 504
rect 6311 391 6345 516
rect 6410 504 6455 515
rect 6421 379 6455 504
rect 6535 379 6569 885
rect 6191 341 6249 379
rect 6283 341 6321 379
rect 6409 341 6467 379
rect 6191 316 6321 341
rect 6373 316 6467 341
rect 6535 375 6557 379
rect 6227 312 6258 316
rect 6398 312 6431 316
rect 6215 307 6299 312
rect 6357 307 6443 312
rect 6225 301 6270 307
rect 6386 301 6433 307
rect 6265 284 6393 293
rect 6253 278 6405 284
rect 6249 273 6409 278
rect 6265 269 6296 273
rect 6360 269 6393 273
rect 6535 259 6569 375
rect 6588 259 6622 1021
rect 6780 959 6818 991
rect 6734 935 6818 959
rect 6827 935 6830 987
rect 6734 919 6890 935
rect 6734 913 6792 919
rect 6748 889 6778 913
rect 6815 889 6890 919
rect 6904 889 6949 1021
rect 6827 885 6858 889
rect 6702 881 6736 885
rect 6790 881 6833 885
rect 6690 851 6748 881
rect 6778 851 6833 881
rect 6904 852 6914 889
rect 6923 885 6949 889
rect 6690 817 6833 851
rect 6923 833 6938 885
rect 6690 779 6748 817
rect 6778 779 6824 817
rect 6904 783 6938 833
rect 6702 693 6736 779
rect 6790 693 6824 779
rect 6793 681 6824 693
rect 6780 677 6824 681
rect 6827 767 6858 783
rect 6780 649 6820 677
rect 6734 609 6820 649
rect 6734 603 6792 609
rect 6807 575 6820 609
rect 6827 655 6861 767
rect 6827 643 6858 655
rect 6827 575 6830 643
rect 6780 569 6818 573
rect 6780 541 6820 569
rect 6734 501 6820 541
rect 6734 495 6792 501
rect 6807 467 6820 501
rect 6827 501 6830 569
rect 6827 489 6858 501
rect 6793 462 6824 467
rect 6691 451 6736 462
rect 6779 451 6824 462
rect 6702 379 6736 451
rect 6790 379 6824 451
rect 6827 391 6861 489
rect 6827 379 6858 391
rect 6690 341 6748 379
rect 6778 375 6858 379
rect 6778 341 6833 375
rect 6690 313 6833 341
rect 6904 341 6949 783
rect 6690 307 6836 313
rect 6690 263 6748 307
rect 6778 263 6836 307
rect 6904 259 6938 341
rect 6957 259 6991 1412
rect 7015 1300 7045 1412
rect 7015 1008 7049 1300
rect 7071 1246 7083 1250
rect 7059 1046 7103 1246
rect 7071 1042 7083 1046
rect 7015 882 7045 1008
rect 7015 590 7049 882
rect 7071 828 7083 832
rect 7059 628 7103 828
rect 7071 624 7083 628
rect 7015 464 7045 590
rect 7015 259 7049 464
rect 7071 410 7083 414
rect 5667 225 6992 259
rect 7034 225 7049 259
rect 7059 225 7103 410
rect 7529 396 7543 2194
rect 7563 442 7597 2194
rect 7651 2140 7663 2160
rect 7751 2142 7797 2173
rect 7669 2140 7709 2142
rect 7651 2126 7709 2140
rect 7739 2127 7797 2142
rect 7719 2126 7797 2127
rect 7651 2081 7797 2126
rect 7851 2093 7863 2099
rect 7851 2081 7881 2093
rect 7895 2081 7929 2194
rect 8291 2175 8306 2209
rect 7663 2077 7691 2081
rect 7751 2077 7785 2081
rect 7623 2045 7657 2049
rect 7781 2045 7815 2049
rect 7611 2043 7657 2045
rect 7741 2043 7815 2045
rect 7611 1845 7651 2043
rect 7741 2034 7791 2043
rect 7707 2000 7791 2034
rect 7747 1994 7753 2000
rect 7775 1966 7791 2000
rect 7909 1984 7929 2081
rect 7741 1896 7788 1909
rect 7741 1862 7791 1896
rect 7914 1878 7929 1984
rect 7707 1845 7791 1862
rect 7623 1841 7631 1845
rect 7707 1832 7741 1836
rect 7747 1832 7757 1845
rect 7781 1841 7791 1845
rect 7691 1828 7793 1832
rect 7695 1822 7707 1828
rect 7741 1822 7753 1828
rect 7673 1803 7707 1804
rect 7741 1803 7765 1804
rect 7673 1798 7765 1803
rect 7663 1790 7789 1798
rect 7663 1781 7709 1790
rect 7739 1781 7789 1790
rect 7909 1781 7929 1878
rect 7654 1766 7797 1781
rect 7669 1764 7797 1766
rect 7669 1748 7709 1764
rect 7739 1748 7769 1764
rect 7651 1690 7663 1724
rect 7751 1706 7797 1737
rect 7669 1690 7709 1706
rect 7739 1690 7797 1706
rect 7669 1656 7797 1690
rect 7669 1647 7709 1656
rect 7623 1609 7657 1613
rect 7611 1543 7657 1609
rect 7663 1609 7709 1647
rect 7739 1627 7785 1656
rect 7739 1609 7815 1627
rect 7663 1593 7697 1609
rect 7751 1593 7815 1609
rect 7663 1577 7691 1593
rect 7611 1409 7651 1543
rect 7781 1421 7815 1593
rect 7851 1581 7881 1663
rect 7895 1581 7929 1781
rect 7909 1484 7929 1581
rect 7623 1405 7631 1409
rect 7914 1379 7929 1484
rect 7669 1312 7769 1350
rect 7651 1270 7697 1288
rect 7751 1282 7787 1288
rect 7909 1282 7929 1379
rect 7751 1270 7797 1282
rect 7651 1254 7663 1270
rect 7669 1254 7709 1270
rect 7739 1254 7797 1270
rect 7669 1220 7797 1254
rect 7669 1211 7709 1220
rect 7623 1173 7657 1177
rect 7611 1044 7657 1173
rect 7663 1173 7709 1211
rect 7739 1173 7785 1220
rect 7663 1094 7697 1173
rect 7751 1161 7785 1173
rect 7751 1094 7815 1161
rect 7663 1078 7691 1094
rect 7781 1082 7815 1094
rect 7851 1082 7881 1227
rect 7895 1082 7929 1282
rect 7611 973 7651 1044
rect 7741 1035 7815 1082
rect 7707 1001 7815 1035
rect 7747 995 7753 1001
rect 7775 985 7815 1001
rect 7909 985 7929 1082
rect 7775 973 7791 985
rect 7623 969 7631 973
rect 7781 969 7791 973
rect 7685 898 7753 902
rect 7669 892 7769 898
rect 7673 886 7707 892
rect 7741 886 7765 892
rect 7914 880 7929 985
rect 7695 864 7707 870
rect 7741 864 7753 870
rect 7691 858 7757 864
rect 7707 852 7741 858
rect 7691 830 7757 852
rect 7663 796 7785 818
rect 7663 787 7669 796
rect 7685 784 7753 796
rect 7769 787 7785 796
rect 7909 783 7929 880
rect 7654 768 7709 783
rect 7623 737 7657 741
rect 7611 545 7657 737
rect 7663 737 7709 768
rect 7739 771 7784 783
rect 7739 737 7785 771
rect 7663 595 7697 737
rect 7751 725 7785 737
rect 7751 595 7815 725
rect 7663 579 7691 595
rect 7781 549 7815 595
rect 7851 583 7881 783
rect 7895 583 7929 783
rect 7816 554 7821 583
rect 7844 582 7849 583
rect 7611 537 7651 545
rect 7623 533 7631 537
rect 7909 502 7929 583
rect 7658 490 7753 498
rect 7658 464 7685 490
rect 7895 464 7929 502
rect 7948 2141 8067 2175
rect 8121 2141 8368 2175
rect 7948 464 7982 2141
rect 8133 2120 8167 2141
rect 8121 2107 8239 2120
rect 8084 2081 8239 2107
rect 8300 2091 8325 2141
rect 8333 2122 8368 2141
rect 8391 2122 8422 2229
rect 8334 2091 8368 2122
rect 8300 2081 8368 2091
rect 8129 2079 8179 2081
rect 8112 2073 8204 2079
rect 8300 2077 8325 2081
rect 8108 2068 8204 2073
rect 8108 2061 8208 2068
rect 8108 2043 8211 2061
rect 8129 2040 8211 2043
rect 8129 2039 8208 2040
rect 8179 2030 8258 2034
rect 8179 2005 8279 2030
rect 8186 2000 8279 2005
rect 8186 1994 8275 2000
rect 8208 1992 8258 1994
rect 8208 1984 8266 1992
rect 8214 1969 8266 1984
rect 8214 1966 8260 1969
rect 8220 1962 8254 1966
rect 8220 1878 8266 1909
rect 8208 1862 8266 1878
rect 8195 1835 8288 1862
rect 8050 1828 8108 1835
rect 8179 1828 8288 1835
rect 8050 1792 8121 1828
rect 8179 1792 8266 1828
rect 8062 1788 8089 1792
rect 8028 1781 8055 1785
rect 8028 1769 8180 1781
rect 8024 1766 8180 1769
rect 8028 1764 8180 1766
rect 8028 1754 8055 1764
rect 8121 1745 8180 1764
rect 8192 1745 8239 1781
rect 8285 1769 8288 1781
rect 8121 1711 8239 1745
rect 8121 1695 8179 1711
rect 8121 1684 8136 1695
rect 8121 1680 8180 1684
rect 8133 1668 8180 1680
rect 8121 1637 8180 1668
rect 8192 1637 8239 1684
rect 7996 1584 8067 1610
rect 8121 1603 8239 1637
rect 8121 1584 8208 1603
rect 7996 1581 8208 1584
rect 8028 1577 8055 1581
rect 8300 1577 8325 1785
rect 8062 1556 8089 1560
rect 8220 1556 8254 1568
rect 8056 1553 8102 1556
rect 8062 1543 8089 1553
rect 8208 1534 8266 1556
rect 8195 1500 8288 1534
rect 8208 1484 8266 1500
rect 8251 1469 8266 1484
rect 8220 1394 8254 1410
rect 8263 1394 8266 1410
rect 8220 1379 8266 1394
rect 8208 1363 8266 1379
rect 8195 1356 8266 1363
rect 8195 1343 8263 1356
rect 8179 1330 8263 1343
rect 8179 1329 8258 1330
rect 8183 1323 8232 1329
rect 8193 1320 8232 1323
rect 8155 1309 8204 1315
rect 8129 1308 8208 1309
rect 8124 1295 8208 1308
rect 8124 1292 8204 1295
rect 8124 1282 8192 1292
rect 8121 1275 8239 1282
rect 8121 1259 8179 1275
rect 8121 1248 8167 1259
rect 8121 1244 8180 1248
rect 8133 1232 8180 1244
rect 8121 1201 8180 1232
rect 8192 1201 8239 1248
rect 8121 1167 8239 1201
rect 8028 1146 8055 1158
rect 8024 1094 8055 1146
rect 8028 1078 8055 1094
rect 8062 1108 8089 1124
rect 8121 1120 8179 1167
rect 8062 1056 8093 1108
rect 8095 1056 8096 1108
rect 8133 1094 8167 1120
rect 8209 1108 8254 1119
rect 8062 1044 8089 1056
rect 8099 1054 8102 1083
rect 8127 1082 8130 1083
rect 8220 1082 8254 1108
rect 8257 1082 8260 1120
rect 8285 1082 8288 1148
rect 8291 1094 8292 1146
rect 8208 1035 8266 1082
rect 8300 1078 8325 1286
rect 8195 1001 8288 1035
rect 8208 985 8266 1001
rect 8251 970 8266 985
rect 8157 839 8192 873
rect 8195 830 8230 864
rect 8133 783 8167 799
rect 8121 765 8180 783
rect 8192 765 8239 783
rect 8121 731 8239 765
rect 8028 710 8055 722
rect 8024 595 8055 710
rect 8028 579 8055 595
rect 8062 672 8089 688
rect 8121 684 8179 731
rect 8062 557 8093 672
rect 8095 557 8096 672
rect 8133 595 8167 684
rect 8209 672 8254 683
rect 8220 583 8254 672
rect 8291 595 8292 710
rect 8062 545 8089 557
rect 8208 536 8266 583
rect 8300 579 8325 787
rect 8050 484 8108 518
rect 8195 502 8288 536
rect 8208 484 8266 502
rect 8062 480 8096 484
rect 8220 480 8254 484
rect 8090 464 8226 471
rect 8334 464 8368 2081
rect 8387 2088 8607 2122
rect 8661 2088 8733 2122
rect 8387 2081 8422 2088
rect 8387 1781 8421 2081
rect 8449 2000 8455 2034
rect 8523 1994 8545 2040
rect 8549 2020 8581 2034
rect 8551 1980 8573 2020
rect 8659 1909 8693 1927
rect 8501 1896 8548 1909
rect 8501 1893 8567 1896
rect 8449 1828 8455 1862
rect 8489 1828 8567 1893
rect 8659 1862 8705 1909
rect 8723 1862 8727 1868
rect 8489 1781 8547 1828
rect 8659 1785 8693 1862
rect 8695 1794 8699 1862
rect 8704 1785 8705 1862
rect 8719 1828 8733 1862
rect 8723 1822 8727 1828
rect 8561 1781 8569 1785
rect 8387 1581 8422 1781
rect 8501 1751 8541 1781
rect 8554 1780 8569 1781
rect 8550 1769 8595 1780
rect 8526 1739 8541 1751
rect 8554 1739 8595 1769
rect 8659 1751 8707 1785
rect 8673 1739 8707 1751
rect 8527 1735 8535 1739
rect 8549 1726 8607 1739
rect 8529 1692 8607 1726
rect 8549 1642 8607 1692
rect 8639 1658 8647 1692
rect 8661 1658 8707 1739
rect 8592 1631 8607 1642
rect 8516 1627 8607 1631
rect 8661 1631 8662 1658
rect 8673 1631 8707 1658
rect 8516 1615 8595 1627
rect 8516 1584 8607 1615
rect 8661 1593 8707 1631
rect 8387 1282 8421 1581
rect 8549 1568 8631 1584
rect 8547 1555 8631 1568
rect 8547 1550 8599 1555
rect 8639 1550 8647 1584
rect 8661 1581 8681 1593
rect 8673 1577 8681 1581
rect 8551 1544 8573 1550
rect 8523 1540 8535 1543
rect 8523 1534 8545 1540
rect 8449 1500 8455 1534
rect 8497 1529 8549 1534
rect 8465 1516 8549 1529
rect 8465 1503 8547 1516
rect 8465 1500 8580 1503
rect 8489 1484 8547 1500
rect 8489 1469 8535 1484
rect 8501 1462 8535 1469
rect 8685 1466 8693 1507
rect 8695 1466 8699 1503
rect 8704 1469 8705 1503
rect 8719 1500 8733 1534
rect 8723 1494 8727 1500
rect 8501 1397 8548 1410
rect 8688 1397 8705 1410
rect 8501 1394 8567 1397
rect 8449 1329 8455 1363
rect 8489 1329 8567 1394
rect 8685 1363 8705 1397
rect 8723 1363 8727 1369
rect 8685 1336 8693 1363
rect 8695 1336 8699 1363
rect 8704 1336 8705 1363
rect 8489 1303 8549 1329
rect 8607 1303 8705 1336
rect 8719 1329 8733 1363
rect 8723 1323 8727 1329
rect 8527 1299 8535 1303
rect 8659 1299 8693 1303
rect 8529 1282 8595 1290
rect 8673 1282 8707 1286
rect 8387 1082 8422 1282
rect 8529 1256 8607 1282
rect 8625 1275 8727 1282
rect 8661 1265 8707 1275
rect 8549 1206 8607 1256
rect 8639 1222 8647 1256
rect 8661 1222 8681 1265
rect 8592 1191 8607 1206
rect 8661 1195 8662 1222
rect 8673 1195 8681 1222
rect 8661 1188 8681 1195
rect 8661 1182 8678 1188
rect 8529 1164 8561 1182
rect 8592 1164 8607 1179
rect 8529 1148 8607 1164
rect 8549 1121 8607 1148
rect 8547 1082 8607 1121
rect 8639 1114 8647 1148
rect 8661 1121 8681 1182
rect 8661 1095 8733 1121
rect 8625 1082 8733 1095
rect 8387 783 8421 1082
rect 8561 1078 8569 1082
rect 8673 1078 8707 1082
rect 8527 1069 8535 1071
rect 8501 1067 8567 1069
rect 8659 1067 8693 1071
rect 8449 1001 8455 1035
rect 8489 1001 8567 1067
rect 8653 1054 8705 1067
rect 8659 1044 8705 1054
rect 8685 1035 8705 1044
rect 8723 1035 8727 1041
rect 8489 985 8547 1001
rect 8489 970 8504 985
rect 8685 967 8693 1035
rect 8695 967 8699 1035
rect 8704 970 8705 1035
rect 8719 1001 8733 1035
rect 8723 995 8727 1001
rect 8489 867 8580 911
rect 8688 898 8705 911
rect 8685 867 8705 898
rect 8497 864 8547 867
rect 8449 830 8455 864
rect 8465 854 8547 864
rect 8685 863 8693 867
rect 8723 864 8727 870
rect 8465 841 8549 854
rect 8497 830 8549 841
rect 8719 830 8733 864
rect 8523 824 8545 830
rect 8551 820 8573 826
rect 8547 809 8599 820
rect 8614 809 8631 820
rect 8547 796 8631 809
rect 8549 786 8631 796
rect 8639 786 8647 820
rect 8549 784 8599 786
rect 8523 783 8599 784
rect 8387 583 8422 783
rect 8549 770 8607 783
rect 8561 755 8607 770
rect 8661 759 8662 783
rect 8673 771 8681 787
rect 8673 759 8707 771
rect 8561 748 8595 755
rect 8529 728 8561 746
rect 8592 728 8607 743
rect 8529 712 8607 728
rect 8527 630 8535 635
rect 8549 631 8607 712
rect 8639 678 8647 712
rect 8661 678 8707 759
rect 8661 631 8662 678
rect 8490 619 8535 630
rect 8501 583 8535 619
rect 8561 595 8595 631
rect 8673 629 8707 678
rect 8659 595 8707 629
rect 8387 464 8421 583
rect 8489 570 8548 583
rect 8561 579 8569 595
rect 8659 583 8693 595
rect 8449 502 8455 536
rect 8489 502 8567 570
rect 8659 536 8705 583
rect 8723 536 8727 542
rect 8489 486 8547 502
rect 8489 471 8535 486
rect 8501 464 8535 471
rect 8659 464 8693 536
rect 8695 468 8699 536
rect 8704 471 8705 536
rect 8719 502 8733 536
rect 8723 496 8727 502
rect 7658 453 8705 464
rect 7669 443 8705 453
rect 7669 442 8733 443
rect 7563 430 8733 442
rect 7914 354 7929 430
rect 7948 354 7982 430
rect 8334 397 8368 430
rect 7948 320 7963 354
rect 8353 301 8368 397
rect 8387 301 8421 430
rect 8467 403 8569 420
rect 8625 403 8727 420
rect 8387 267 8402 301
rect 5686 195 5974 225
rect 6055 195 6070 225
rect 6089 195 6123 225
rect 5314 172 5372 178
rect 5314 138 5326 172
rect 6089 161 6104 195
rect 6554 142 6569 224
rect 6588 142 6622 225
rect 6734 191 6746 225
rect 6734 185 6792 191
rect 6904 185 6938 225
rect 5314 132 5372 138
rect 6588 108 6603 142
rect 6923 89 6938 185
rect 6957 89 6991 225
rect 7071 206 7083 225
rect 3299 55 3314 89
rect 5168 55 5183 89
rect 6957 55 6972 89
<< error_ps >>
rect 8733 2088 8807 2122
rect 8773 1984 8807 2088
rect 8773 1484 8807 1878
rect 8773 985 8807 1379
rect 8826 1163 8877 1197
rect 8931 1163 9077 1197
rect 8826 1082 8860 1163
rect 8986 1082 8989 1111
rect 9019 1095 9077 1111
rect 9002 1082 9077 1095
rect 8773 486 8807 880
rect 8971 985 8986 1014
rect 8987 1001 9021 1014
rect 8971 814 8986 880
rect 8987 830 9021 864
rect 9131 814 9144 1014
rect 8826 583 8860 783
rect 8986 717 8989 783
rect 9019 767 9077 783
rect 9002 733 9077 767
rect 9019 717 9077 733
rect 8986 583 8989 675
rect 9019 659 9077 675
rect 9002 625 9077 659
rect 9019 583 9077 625
rect 9131 464 9144 578
rect 8928 430 9144 464
use pmos_cs  x1
timestamp 1729443144
transform 1 0 254 0 1 1247
box -254 -1247 3431 2093
use pmos_out2  x2
timestamp 1729443144
transform 1 0 7815 0 1 1981
box -342 -1981 2644 500
use nmosdp  x3
timestamp 1729443144
transform 1 0 4031 0 1 799
box -346 -799 1523 798
use nmoscs2  x4
timestamp 1729443144
transform 1 0 5783 0 1 801
box -229 -801 1690 1232
<< end >>
