magic
tech sky130A
magscale 1 2
timestamp 1729443144
<< error_p >>
rect -29 835 29 841
rect -29 801 -17 835
rect -29 795 29 801
rect -29 507 29 513
rect -29 473 -17 507
rect -29 467 29 473
rect -29 399 29 405
rect -29 365 -17 399
rect -29 359 29 365
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect -29 -405 29 -399
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect -29 -513 29 -507
rect -29 -801 29 -795
rect -29 -835 -17 -801
rect -29 -841 29 -835
<< nwell >>
rect -211 -973 211 973
<< pmos >>
rect -15 554 15 754
rect -15 118 15 318
rect -15 -318 15 -118
rect -15 -754 15 -554
<< pdiff >>
rect -73 742 -15 754
rect -73 566 -61 742
rect -27 566 -15 742
rect -73 554 -15 566
rect 15 742 73 754
rect 15 566 27 742
rect 61 566 73 742
rect 15 554 73 566
rect -73 306 -15 318
rect -73 130 -61 306
rect -27 130 -15 306
rect -73 118 -15 130
rect 15 306 73 318
rect 15 130 27 306
rect 61 130 73 306
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -306 -61 -130
rect -27 -306 -15 -130
rect -73 -318 -15 -306
rect 15 -130 73 -118
rect 15 -306 27 -130
rect 61 -306 73 -130
rect 15 -318 73 -306
rect -73 -566 -15 -554
rect -73 -742 -61 -566
rect -27 -742 -15 -566
rect -73 -754 -15 -742
rect 15 -566 73 -554
rect 15 -742 27 -566
rect 61 -742 73 -566
rect 15 -754 73 -742
<< pdiffc >>
rect -61 566 -27 742
rect 27 566 61 742
rect -61 130 -27 306
rect 27 130 61 306
rect -61 -306 -27 -130
rect 27 -306 61 -130
rect -61 -742 -27 -566
rect 27 -742 61 -566
<< nsubdiff >>
rect -175 903 -79 937
rect 79 903 175 937
rect -175 841 -141 903
rect 141 841 175 903
rect -175 -903 -141 -841
rect 141 -903 175 -841
rect -175 -937 -79 -903
rect 79 -937 175 -903
<< nsubdiffcont >>
rect -79 903 79 937
rect -175 -841 -141 841
rect 141 -841 175 841
rect -79 -937 79 -903
<< poly >>
rect -33 835 33 851
rect -33 801 -17 835
rect 17 801 33 835
rect -33 785 33 801
rect -15 754 15 785
rect -15 523 15 554
rect -33 507 33 523
rect -33 473 -17 507
rect 17 473 33 507
rect -33 457 33 473
rect -33 399 33 415
rect -33 365 -17 399
rect 17 365 33 399
rect -33 349 33 365
rect -15 318 15 349
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -349 15 -318
rect -33 -365 33 -349
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -415 33 -399
rect -33 -473 33 -457
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -33 -523 33 -507
rect -15 -554 15 -523
rect -15 -785 15 -754
rect -33 -801 33 -785
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -33 -851 33 -835
<< polycont >>
rect -17 801 17 835
rect -17 473 17 507
rect -17 365 17 399
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -17 -835 17 -801
<< locali >>
rect -175 903 -79 937
rect 79 903 175 937
rect -175 841 -141 903
rect 141 841 175 903
rect -33 801 -17 835
rect 17 801 33 835
rect -61 742 -27 758
rect -61 550 -27 566
rect 27 742 61 758
rect 27 550 61 566
rect -33 473 -17 507
rect 17 473 33 507
rect -33 365 -17 399
rect 17 365 33 399
rect -61 306 -27 322
rect -61 114 -27 130
rect 27 306 61 322
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -322 -27 -306
rect 27 -130 61 -114
rect 27 -322 61 -306
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -507 -17 -473
rect 17 -507 33 -473
rect -61 -566 -27 -550
rect -61 -758 -27 -742
rect 27 -566 61 -550
rect 27 -758 61 -742
rect -33 -835 -17 -801
rect 17 -835 33 -801
rect -175 -903 -141 -841
rect 141 -903 175 -841
rect -175 -937 -79 -903
rect 79 -937 175 -903
<< viali >>
rect -17 801 17 835
rect -61 566 -27 742
rect 27 566 61 742
rect -17 473 17 507
rect -17 365 17 399
rect -61 130 -27 306
rect 27 130 61 306
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -306 -27 -130
rect 27 -306 61 -130
rect -17 -399 17 -365
rect -17 -507 17 -473
rect -61 -742 -27 -566
rect 27 -742 61 -566
rect -17 -835 17 -801
<< metal1 >>
rect -29 835 29 841
rect -29 801 -17 835
rect 17 801 29 835
rect -29 795 29 801
rect -67 742 -21 754
rect -67 566 -61 742
rect -27 566 -21 742
rect -67 554 -21 566
rect 21 742 67 754
rect 21 566 27 742
rect 61 566 67 742
rect 21 554 67 566
rect -29 507 29 513
rect -29 473 -17 507
rect 17 473 29 507
rect -29 467 29 473
rect -29 399 29 405
rect -29 365 -17 399
rect 17 365 29 399
rect -29 359 29 365
rect -67 306 -21 318
rect -67 130 -61 306
rect -27 130 -21 306
rect -67 118 -21 130
rect 21 306 67 318
rect 21 130 27 306
rect 61 130 67 306
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -306 -61 -130
rect -27 -306 -21 -130
rect -67 -318 -21 -306
rect 21 -130 67 -118
rect 21 -306 27 -130
rect 61 -306 67 -130
rect 21 -318 67 -306
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect 17 -399 29 -365
rect -29 -405 29 -399
rect -29 -473 29 -467
rect -29 -507 -17 -473
rect 17 -507 29 -473
rect -29 -513 29 -507
rect -67 -566 -21 -554
rect -67 -742 -61 -566
rect -27 -742 -21 -566
rect -67 -754 -21 -742
rect 21 -566 67 -554
rect 21 -742 27 -566
rect 61 -742 67 -566
rect 21 -754 67 -742
rect -29 -801 29 -795
rect -29 -835 -17 -801
rect 17 -835 29 -801
rect -29 -841 29 -835
<< properties >>
string FIXED_BBOX -158 -920 158 920
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
