magic
tech sky130A
magscale 1 2
timestamp 1729440139
<< checkpaint >>
rect 690 835 3632 888
rect 690 -3578 4001 835
rect 1059 -3631 4001 -3578
<< error_s >>
rect 3 205 26 228
rect 54 205 77 228
rect 105 214 228 228
rect 161 205 228 214
rect 0 177 26 200
rect 54 186 200 200
rect 54 177 105 186
rect 133 177 200 186
rect 0 0 12 20
rect 68 0 170 20
rect -28 -20 -16 -8
rect -22 -28 -16 -20
rect 96 -28 142 -8
rect -156 -177 211 -143
rect -181 -208 -175 -177
rect -156 -208 -121 -177
rect -91 -198 -68 -187
rect -56 -198 -16 -177
rect -91 -208 82 -198
rect -178 -239 -175 -208
rect -144 -212 -141 -208
rect -91 -229 -68 -208
rect -56 -212 -22 -208
rect -49 -234 -26 -229
rect 0 -236 12 -208
rect -49 -246 35 -245
rect 0 -249 35 -246
rect 0 -255 49 -249
rect 0 -279 74 -255
rect 6 -288 74 -279
rect 6 -289 90 -288
rect 148 -289 164 -255
rect 177 -305 211 -177
rect 576 -196 588 -162
rect 664 -195 684 -162
rect 652 -196 710 -195
rect 177 -316 188 -305
rect 63 -323 97 -322
rect 0 -400 57 -393
rect 63 -411 109 -380
rect 196 -393 211 -305
rect 133 -400 211 -393
rect 51 -421 109 -411
rect 177 -411 188 -400
rect 196 -411 211 -400
rect 177 -421 211 -411
rect 230 -208 710 -196
rect 230 -217 248 -208
rect 306 -217 406 -208
rect 464 -217 564 -208
rect 230 -230 270 -217
rect 284 -221 428 -217
rect 442 -221 586 -217
rect 272 -230 598 -221
rect 615 -230 650 -208
rect 664 -212 684 -208
rect 230 -289 264 -230
rect 616 -249 650 -230
rect 306 -264 406 -255
rect 356 -275 406 -264
rect 464 -264 564 -255
rect 464 -267 524 -264
rect 356 -282 420 -275
rect 356 -289 406 -282
rect 458 -289 524 -267
rect 230 -305 248 -289
rect 366 -295 393 -289
rect 458 -292 477 -289
rect 394 -298 421 -292
rect 230 -411 264 -305
rect 390 -323 490 -298
rect 406 -327 419 -323
rect 451 -327 474 -323
rect 344 -396 437 -380
rect 3 -428 109 -421
rect 161 -427 228 -421
rect -209 -508 -175 -454
rect 6 -461 109 -428
rect 148 -428 223 -427
rect 148 -461 164 -428
rect 51 -470 90 -461
rect -95 -480 -61 -470
rect -144 -508 -141 -504
rect -129 -508 -110 -504
rect -181 -708 -175 -508
rect -156 -554 -104 -508
rect -101 -526 -61 -480
rect -55 -504 -34 -498
rect -95 -530 -61 -526
rect -56 -509 -27 -504
rect 51 -508 97 -470
rect 103 -504 124 -498
rect -56 -526 -22 -509
rect 63 -514 97 -508
rect 68 -526 97 -514
rect -56 -539 -10 -526
rect -156 -564 -110 -554
rect -67 -564 -10 -539
rect -156 -708 -121 -564
rect -67 -573 -56 -564
rect -49 -573 -10 -564
rect 35 -530 97 -526
rect 102 -520 131 -504
rect 35 -573 82 -530
rect 102 -552 135 -520
rect 102 -564 131 -552
rect -49 -607 82 -573
rect -49 -623 -10 -607
rect -67 -649 -56 -647
rect -28 -649 -16 -623
rect -80 -662 -16 -649
rect 0 -662 12 -613
rect -80 -675 12 -662
rect -80 -681 0 -675
rect 35 -681 82 -634
rect -80 -696 82 -681
rect -64 -708 82 -696
rect -178 -746 -175 -708
rect -144 -712 -141 -708
rect -49 -715 -10 -708
rect -49 -734 -26 -715
rect 29 -755 74 -740
rect 51 -762 97 -755
rect 6 -789 109 -762
rect 148 -789 164 -755
rect 51 -805 90 -789
rect 177 -805 211 -428
rect 177 -816 188 -805
rect 29 -911 53 -872
rect 57 -880 81 -872
rect 57 -911 109 -880
rect 29 -921 109 -911
rect 31 -927 109 -921
rect 177 -911 188 -900
rect 196 -911 211 -805
rect 6 -930 109 -927
rect -49 -954 -26 -940
rect 6 -954 131 -930
rect -209 -1008 -175 -954
rect -107 -962 -26 -954
rect -10 -962 131 -954
rect 148 -961 164 -927
rect -49 -986 -26 -962
rect -144 -1008 -141 -1004
rect -49 -1008 12 -986
rect 105 -990 131 -962
rect -181 -1208 -175 -1008
rect -156 -1160 -121 -1008
rect -80 -1009 12 -1008
rect 35 -1009 82 -1008
rect -64 -1023 82 -1009
rect -49 -1043 82 -1023
rect -49 -1059 -10 -1043
rect -67 -1117 -56 -1083
rect -28 -1101 -16 -1059
rect -49 -1117 -10 -1101
rect 0 -1111 12 -1049
rect 35 -1117 82 -1070
rect -49 -1151 82 -1117
rect -49 -1160 -10 -1151
rect -156 -1170 -110 -1160
rect -156 -1208 -104 -1170
rect -83 -1194 -62 -1180
rect -95 -1198 -61 -1194
rect -178 -1246 -175 -1208
rect -144 -1212 -141 -1208
rect -129 -1212 -110 -1208
rect -101 -1236 -61 -1198
rect -56 -1198 -10 -1160
rect -56 -1208 -16 -1198
rect 0 -1200 12 -1157
rect 102 -1172 131 -1160
rect 68 -1199 97 -1194
rect 52 -1208 97 -1199
rect -56 -1212 -27 -1208
rect 51 -1210 97 -1208
rect 102 -1196 135 -1172
rect 102 -1210 131 -1196
rect 51 -1212 131 -1210
rect -95 -1246 -61 -1236
rect 51 -1255 109 -1212
rect 6 -1289 109 -1255
rect 148 -1289 164 -1255
rect 51 -1305 90 -1289
rect 177 -1305 211 -911
rect 177 -1316 188 -1305
rect 57 -1398 103 -1372
rect 29 -1426 131 -1400
rect 196 -2017 211 -1305
rect 230 -508 248 -411
rect 252 -508 264 -454
rect 332 -461 437 -396
rect 502 -411 548 -380
rect 490 -427 548 -411
rect 480 -461 570 -427
rect 332 -508 390 -461
rect 490 -508 548 -461
rect 635 -470 650 -249
rect 230 -708 264 -508
rect 344 -567 378 -508
rect 407 -520 452 -509
rect 418 -579 452 -520
rect 502 -567 536 -508
rect 406 -626 465 -579
rect 474 -626 521 -579
rect 406 -660 521 -626
rect 406 -676 464 -660
rect 359 -708 521 -687
rect 230 -805 248 -708
rect 418 -712 452 -708
rect 582 -712 610 -504
rect 394 -734 486 -728
rect 372 -746 486 -734
rect 372 -749 390 -746
rect 366 -768 393 -749
rect 322 -777 393 -768
rect 394 -768 424 -746
rect 446 -755 474 -746
rect 490 -755 498 -734
rect 616 -746 650 -470
rect 669 -283 704 -249
rect 669 -504 703 -283
rect 1186 -344 1379 41
rect 1696 -343 2050 -118
rect 1696 -344 1762 -343
rect 664 -708 703 -504
rect 2132 -510 2190 -504
rect 2132 -544 2144 -510
rect 2132 -550 2190 -544
rect 664 -712 684 -708
rect 451 -768 474 -755
rect 480 -768 512 -755
rect 394 -774 421 -768
rect 480 -777 548 -768
rect 310 -789 406 -777
rect 468 -789 564 -777
rect 319 -795 342 -789
rect 366 -795 393 -789
rect 477 -795 551 -789
rect 478 -798 550 -795
rect 230 -911 264 -805
rect 344 -815 378 -811
rect 502 -815 536 -811
rect 332 -820 390 -815
rect 490 -820 548 -815
rect 338 -823 342 -820
rect 344 -823 384 -820
rect 496 -826 542 -820
rect 344 -896 437 -880
rect 230 -1008 248 -911
rect 252 -1008 264 -954
rect 332 -961 437 -896
rect 502 -911 548 -880
rect 490 -927 548 -911
rect 480 -961 570 -927
rect 332 -1008 390 -961
rect 490 -1008 548 -961
rect 635 -970 650 -746
rect 230 -1208 264 -1008
rect 407 -1015 452 -1009
rect 406 -1062 465 -1015
rect 474 -1062 521 -1015
rect 406 -1096 521 -1062
rect 406 -1112 464 -1096
rect 418 -1154 465 -1123
rect 406 -1170 465 -1154
rect 474 -1170 521 -1123
rect 406 -1197 521 -1170
rect 390 -1204 521 -1197
rect 390 -1208 490 -1204
rect 230 -1305 248 -1208
rect 582 -1212 610 -1004
rect 310 -1251 412 -1229
rect 310 -1255 437 -1251
rect 310 -1263 322 -1255
rect 332 -1289 437 -1255
rect 468 -1263 570 -1229
rect 616 -1246 650 -970
rect 669 -734 684 -712
rect 669 -1004 703 -734
rect 2132 -838 2190 -832
rect 2132 -872 2144 -838
rect 2132 -878 2190 -872
rect 2132 -946 2190 -940
rect 2132 -980 2144 -946
rect 2132 -986 2190 -980
rect 664 -1208 703 -1004
rect 1055 -1174 1089 -1120
rect 664 -1212 684 -1208
rect 480 -1289 570 -1263
rect 332 -1305 390 -1289
rect 490 -1305 548 -1289
rect 230 -2017 264 -1305
rect 332 -1320 347 -1305
rect 533 -1320 548 -1305
rect 230 -2051 245 -2017
rect 635 -2070 650 -1246
rect 669 -1234 684 -1212
rect 669 -2070 703 -1234
rect 669 -2104 684 -2070
rect 1074 -2123 1089 -1174
rect 1108 -1208 1143 -1174
rect 1493 -1208 1528 -1174
rect 1108 -2123 1142 -1208
rect 1494 -1227 1528 -1208
rect 1108 -2157 1123 -2123
rect 1513 -2176 1528 -1227
rect 1547 -1261 1582 -1227
rect 1547 -2176 1581 -1261
rect 1547 -2210 1562 -2176
rect 1952 -2229 1967 -1227
rect 1986 -2229 2020 -1173
rect 2132 -1274 2190 -1268
rect 2132 -1308 2144 -1274
rect 2132 -1314 2190 -1308
rect 2132 -1382 2190 -1376
rect 2132 -1416 2144 -1382
rect 2132 -1422 2190 -1416
rect 2132 -1710 2190 -1704
rect 2132 -1744 2144 -1710
rect 2132 -1750 2190 -1744
rect 2132 -1818 2190 -1812
rect 2132 -1852 2144 -1818
rect 2132 -1858 2190 -1852
rect 2132 -2146 2190 -2140
rect 2132 -2180 2144 -2146
rect 2132 -2186 2190 -2180
rect 1986 -2263 2001 -2229
<< nwell >>
rect -192 -289 746 592
rect -192 -307 184 -289
rect 212 -306 342 -289
rect 370 -306 746 -289
rect 212 -307 746 -306
rect -192 -1308 746 -307
<< poly >>
rect 464 -289 564 -288
rect 15 -461 67 -460
<< metal1 >>
rect 263 304 291 308
rect 105 242 133 304
rect 260 292 294 304
rect 263 242 291 292
rect 421 242 449 304
rect 26 200 54 225
rect 105 214 449 242
rect 0 156 200 200
rect 0 54 212 156
rect 0 0 200 54
rect 0 -400 200 -200
rect 184 -427 212 -426
rect 0 -789 200 -600
rect 0 -800 212 -789
rect 184 -844 212 -800
rect 25 -872 212 -844
rect 25 -927 53 -872
rect 263 -930 291 214
rect 499 156 527 211
rect 341 128 527 156
rect 341 73 369 128
rect 342 -427 370 -425
rect 342 -844 370 -789
rect 478 -798 550 -746
rect 342 -872 528 -844
rect 500 -927 528 -872
rect 105 -958 449 -930
rect 105 -1000 133 -958
rect 0 -1200 200 -1000
rect 263 -1031 291 -958
rect 421 -1021 449 -958
rect 266 -1207 288 -1031
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729312887
transform 1 0 637 0 1 -1108
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729312887
transform 1 0 -83 0 1 392
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729312887
transform 1 0 -83 0 1 -108
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729312887
transform 1 0 637 0 1 -108
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729312887
transform 1 0 -83 0 1 -608
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729312887
transform 1 0 637 0 1 -608
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729312887
transform 1 0 -83 0 1 -1108
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_8
timestamp 1729312887
transform 1 0 637 0 1 392
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHRSS5  sky130_fd_pr__pfet_01v8_BHRSS5_1
timestamp 1729334953
transform 1 0 1330 0 1 -144
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_BHRSS5  sky130_fd_pr__pfet_01v8_BHRSS5_2
timestamp 1729334953
transform 1 0 1618 0 1 -144
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_BHRSS5  sky130_fd_pr__pfet_01v8_BHRSS5_3
timestamp 1729334953
transform 1 0 1906 0 1 -143
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_BHRSS5  sky130_fd_pr__pfet_01v8_BHRSS5_4
timestamp 1729334953
transform 1 0 1906 0 1 -143
box -144 -200 144 200
use sky130_fd_pr__pfet_01v8_V8EU5L  sky130_fd_pr__pfet_01v8_V8EU5L_0
timestamp 1729192300
transform 1 0 277 0 1 392
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_V8EU5L  sky130_fd_pr__pfet_01v8_V8EU5L_1
timestamp 1729192300
transform 1 0 277 0 1 -1108
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_V8EU5L  sky130_fd_pr__pfet_01v8_V8EU5L_2
timestamp 1729192300
transform 1 0 277 0 1 -608
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_V8EU5L  sky130_fd_pr__pfet_01v8_V8EU5L_3
timestamp 1729192300
transform 1 0 277 0 1 -108
box -381 -200 381 200
use sky130_fd_pr__pfet_01v8_XPY429  XM1
timestamp 0
transform 1 0 879 0 1 -1186
box -246 -973 246 973
use sky130_fd_pr__pfet_01v8_XPYQY6  XM2
timestamp 0
transform 1 0 1318 0 1 -1675
box -246 -537 246 537
use sky130_fd_pr__pfet_01v8_XPYQY6  XM3
timestamp 0
transform 1 0 1757 0 1 -1728
box -246 -537 246 537
use sky130_fd_pr__pfet_01v8_XGS9DL  XM4
timestamp 0
transform 1 0 2161 0 1 -1345
box -211 -973 211 973
use sky130_fd_pr__pfet_01v8_XGS9DL  XM5
timestamp 0
transform 1 0 2530 0 1 -1398
box -211 -973 211 973
use sky130_fd_pr__pfet_01v8_XPY429  XM6
timestamp 0
transform 1 0 1 0 1 -1080
box -246 -973 246 973
use sky130_fd_pr__pfet_01v8_XPY429  XM7
timestamp 0
transform 1 0 440 0 1 -1133
box -246 -973 246 973
<< labels >>
flabel nwell 263 -1031 291 308 0 FreeSans 800 0 0 0 S
flabel nwell 464 245 564 292 0 FreeSans 800 0 0 0 M7
flabel nwell -10 245 90 292 0 FreeSans 800 0 0 0 M6
flabel nwell 569 288 705 496 0 FreeSans 800 0 0 0 D7
flabel nwell -151 293 -15 501 0 FreeSans 800 0 0 0 D6
flabel nwell 564 -1212 700 -1004 0 FreeSans 800 0 0 0 D6
flabel nwell -158 -1209 -22 -1001 0 FreeSans 800 0 0 0 D7
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 D5
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VIP
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 OUT
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 D8
port 5 nsew
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
