magic
tech sky130A
magscale 1 2
timestamp 1729443144
<< error_p >>
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect -29 -587 29 -581
<< pwell >>
rect -211 -719 211 719
<< nmos >>
rect -15 109 15 509
rect -15 -509 15 -109
<< ndiff >>
rect -73 497 -15 509
rect -73 121 -61 497
rect -27 121 -15 497
rect -73 109 -15 121
rect 15 497 73 509
rect 15 121 27 497
rect 61 121 73 497
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -497 -61 -121
rect -27 -497 -15 -121
rect -73 -509 -15 -497
rect 15 -121 73 -109
rect 15 -497 27 -121
rect 61 -497 73 -121
rect 15 -509 73 -497
<< ndiffc >>
rect -61 121 -27 497
rect 27 121 61 497
rect -61 -497 -27 -121
rect 27 -497 61 -121
<< psubdiff >>
rect -175 649 -79 683
rect 79 649 175 683
rect -175 587 -141 649
rect 141 587 175 649
rect -175 -649 -141 -587
rect 141 -649 175 -587
rect -175 -683 -79 -649
rect 79 -683 175 -649
<< psubdiffcont >>
rect -79 649 79 683
rect -175 -587 -141 587
rect 141 -587 175 587
rect -79 -683 79 -649
<< poly >>
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -15 509 15 531
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -531 15 -509
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
<< polycont >>
rect -17 547 17 581
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -581 17 -547
<< locali >>
rect -175 649 -79 683
rect 79 649 175 683
rect -175 587 -141 649
rect 141 587 175 649
rect -33 547 -17 581
rect 17 547 33 581
rect -61 497 -27 513
rect -61 105 -27 121
rect 27 497 61 513
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -513 -27 -497
rect 27 -121 61 -105
rect 27 -513 61 -497
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -175 -649 -141 -587
rect 141 -649 175 -587
rect -175 -683 -79 -649
rect 79 -683 175 -649
<< viali >>
rect -17 547 17 581
rect -61 121 -27 497
rect 27 121 61 497
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -497 -27 -121
rect 27 -497 61 -121
rect -17 -581 17 -547
<< metal1 >>
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -67 497 -21 509
rect -67 121 -61 497
rect -27 121 -21 497
rect -67 109 -21 121
rect 21 497 67 509
rect 21 121 27 497
rect 61 121 67 497
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -497 -61 -121
rect -27 -497 -21 -121
rect -67 -509 -21 -497
rect 21 -121 67 -109
rect 21 -497 27 -121
rect 61 -497 67 -121
rect 21 -509 67 -497
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
<< properties >>
string FIXED_BBOX -158 -666 158 666
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
