magic
tech sky130A
magscale 1 2
timestamp 1729443144
<< error_p >>
rect -29 599 29 605
rect -29 565 -17 599
rect -29 559 29 565
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect -29 -605 29 -599
<< nwell >>
rect -211 -737 211 737
<< pmos >>
rect -15 118 15 518
rect -15 -518 15 -118
<< pdiff >>
rect -73 506 -15 518
rect -73 130 -61 506
rect -27 130 -15 506
rect -73 118 -15 130
rect 15 506 73 518
rect 15 130 27 506
rect 61 130 73 506
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -506 -61 -130
rect -27 -506 -15 -130
rect -73 -518 -15 -506
rect 15 -130 73 -118
rect 15 -506 27 -130
rect 61 -506 73 -130
rect 15 -518 73 -506
<< pdiffc >>
rect -61 130 -27 506
rect 27 130 61 506
rect -61 -506 -27 -130
rect 27 -506 61 -130
<< nsubdiff >>
rect -175 667 -79 701
rect 79 667 175 701
rect -175 605 -141 667
rect 141 605 175 667
rect -175 -667 -141 -605
rect 141 -667 175 -605
rect -175 -701 -79 -667
rect 79 -701 175 -667
<< nsubdiffcont >>
rect -79 667 79 701
rect -175 -605 -141 605
rect 141 -605 175 605
rect -79 -701 79 -667
<< poly >>
rect -33 599 33 615
rect -33 565 -17 599
rect 17 565 33 599
rect -33 549 33 565
rect -15 518 15 549
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -549 15 -518
rect -33 -565 33 -549
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -33 -615 33 -599
<< polycont >>
rect -17 565 17 599
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -599 17 -565
<< locali >>
rect -175 667 -79 701
rect 79 667 175 701
rect -175 605 -141 667
rect 141 605 175 667
rect -33 565 -17 599
rect 17 565 33 599
rect -61 506 -27 522
rect -61 114 -27 130
rect 27 506 61 522
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -522 -27 -506
rect 27 -130 61 -114
rect 27 -522 61 -506
rect -33 -599 -17 -565
rect 17 -599 33 -565
rect -175 -667 -141 -605
rect 141 -667 175 -605
rect -175 -701 -79 -667
rect 79 -701 175 -667
<< viali >>
rect -17 565 17 599
rect -61 130 -27 506
rect 27 130 61 506
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -506 -27 -130
rect 27 -506 61 -130
rect -17 -599 17 -565
<< metal1 >>
rect -29 599 29 605
rect -29 565 -17 599
rect 17 565 29 599
rect -29 559 29 565
rect -67 506 -21 518
rect -67 130 -61 506
rect -27 130 -21 506
rect -67 118 -21 130
rect 21 506 67 518
rect 21 130 27 506
rect 61 130 67 506
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -506 -61 -130
rect -27 -506 -21 -130
rect -67 -518 -21 -506
rect 21 -130 67 -118
rect 21 -506 27 -130
rect 61 -506 67 -130
rect 21 -518 67 -506
rect -29 -565 29 -559
rect -29 -599 -17 -565
rect 17 -599 29 -565
rect -29 -605 29 -599
<< properties >>
string FIXED_BBOX -158 -684 158 684
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
