magic
tech sky130A
magscale 1 2
timestamp 1729443867
<< nwell >>
rect -201 1185 834 2093
rect -201 1184 0 1185
rect 81 1184 834 1185
rect -201 -616 834 1184
rect -201 -712 604 -616
rect 696 -665 834 -616
rect 633 -712 834 -665
rect -201 -823 834 -712
<< nsubdiff >>
rect -165 2023 -105 2057
rect 738 2023 798 2057
rect -165 1997 -131 2023
rect 764 1997 798 2023
rect -165 -753 -131 -727
rect 764 -753 798 -727
rect -165 -787 -105 -753
rect 738 -787 798 -753
<< nsubdiffcont >>
rect -105 2023 738 2057
rect -165 -727 -131 1997
rect 764 -727 798 1997
rect -105 -787 738 -753
<< poly >>
rect -62 1973 30 1988
rect -62 1939 -46 1973
rect -12 1939 30 1973
rect -62 1924 30 1939
rect 0 1910 30 1924
rect 604 1966 696 1981
rect 604 1932 646 1966
rect 680 1932 696 1966
rect 604 1917 696 1932
rect 604 1909 634 1917
rect -62 1265 30 1280
rect 88 1272 288 1395
rect -62 1231 -46 1265
rect -12 1231 30 1265
rect -62 1216 30 1231
rect 0 1184 30 1216
rect 604 1265 696 1280
rect 604 1231 646 1265
rect 680 1231 696 1265
rect 604 1216 696 1231
rect 604 1184 634 1216
rect 88 565 546 703
rect 0 52 30 72
rect -62 37 30 52
rect -62 3 -46 37
rect -12 3 30 37
rect -62 -12 30 3
rect 604 51 634 83
rect 604 36 696 51
rect 604 2 646 36
rect 680 2 696 36
rect 346 -128 546 -4
rect 604 -13 696 2
rect 0 -648 30 -629
rect -62 -663 30 -648
rect -62 -697 -46 -663
rect -12 -697 30 -663
rect -62 -712 30 -697
rect 604 -648 634 -628
rect 604 -663 696 -648
rect 604 -697 646 -663
rect 680 -697 696 -663
rect 604 -712 696 -697
<< polycont >>
rect -46 1939 -12 1973
rect 646 1932 680 1966
rect -46 1231 -12 1265
rect 646 1231 680 1265
rect -46 3 -12 37
rect 646 2 680 36
rect -46 -697 -12 -663
rect 646 -697 680 -663
<< locali >>
rect -165 2023 -105 2057
rect 738 2023 798 2057
rect -165 1997 -131 2023
rect 764 1997 798 2023
rect -62 1939 -46 1973
rect -12 1939 4 1973
rect -46 1880 -12 1939
rect 630 1932 646 1966
rect 680 1932 696 1966
rect 646 1868 680 1932
rect -62 1231 -46 1265
rect -12 1231 4 1265
rect 630 1231 646 1265
rect 680 1231 696 1265
rect -46 1184 -12 1231
rect 646 1184 680 1231
rect -46 37 -12 84
rect -62 3 -46 37
rect -12 3 4 37
rect 646 36 680 83
rect 630 2 646 36
rect 680 2 696 36
rect -46 -663 -12 -595
rect 646 -663 680 -601
rect -62 -697 -46 -663
rect -12 -697 4 -663
rect 630 -697 646 -663
rect 680 -697 696 -663
rect -165 -753 -131 -727
rect 764 -753 798 -727
rect -165 -787 -105 -753
rect 738 -787 798 -753
<< viali >>
rect 646 2023 680 2057
rect -46 1939 -12 1973
rect 646 1932 680 1966
rect -46 1231 -12 1265
rect 646 1231 680 1265
rect -46 3 -12 37
rect 646 2 680 36
rect -46 -697 -12 -663
rect 646 -697 680 -663
rect -46 -787 -12 -753
<< metal1 >>
rect 634 2057 692 2063
rect 634 2023 646 2057
rect 680 2023 692 2057
rect -62 1973 0 1979
rect -62 1939 -46 1973
rect -12 1939 0 1973
rect -62 1933 0 1939
rect 634 1972 692 2023
rect 634 1966 696 1972
rect -62 1924 -6 1933
rect 634 1932 646 1966
rect 680 1932 696 1966
rect 634 1926 696 1932
rect -51 1884 -6 1924
rect 640 1917 696 1926
rect 640 1884 685 1917
rect -52 1882 81 1884
rect -56 1872 81 1882
rect -2 1496 81 1872
rect -56 1484 81 1496
rect 300 1435 334 1879
rect 552 1485 685 1884
rect 552 1484 684 1485
rect 604 1435 634 1484
rect 300 1405 634 1435
rect -62 1265 0 1271
rect -62 1231 -46 1265
rect -12 1231 0 1265
rect -62 1216 0 1231
rect -52 1184 0 1216
rect -52 1165 81 1184
rect -51 844 81 1165
rect -51 784 33 844
rect 85 784 95 844
rect -6 527 135 569
rect -6 484 36 527
rect -52 210 82 484
rect -52 84 83 210
rect -52 52 -6 84
rect -62 43 -6 52
rect -62 37 0 43
rect -62 3 -46 37
rect -12 3 0 37
rect -62 -3 0 3
rect 300 -137 334 1405
rect 634 1265 696 1271
rect 634 1231 646 1265
rect 680 1231 696 1265
rect 634 1225 696 1231
rect 640 1216 696 1225
rect 640 1184 685 1216
rect 552 784 685 1184
rect 598 741 640 784
rect 499 699 640 741
rect 539 424 549 484
rect 601 424 686 484
rect 552 84 686 424
rect 634 52 686 84
rect 634 51 692 52
rect 634 36 696 51
rect 634 2 646 36
rect 680 2 696 36
rect 634 -4 696 2
rect 0 -167 334 -137
rect 0 -216 30 -167
rect -52 -594 81 -216
rect -51 -615 81 -594
rect 300 -611 334 -167
rect 552 -228 692 -216
rect 552 -604 638 -228
rect 552 -613 692 -604
rect -51 -648 -6 -615
rect 552 -616 685 -613
rect -62 -657 -6 -648
rect 640 -648 685 -616
rect 640 -657 696 -648
rect -62 -663 0 -657
rect -62 -697 -46 -663
rect -12 -697 0 -663
rect -62 -703 0 -697
rect 634 -663 696 -657
rect 634 -697 646 -663
rect 680 -697 696 -663
rect 634 -703 696 -697
rect -58 -753 0 -703
rect -58 -787 -46 -753
rect -12 -787 0 -753
rect -58 -793 0 -787
<< via1 >>
rect -56 1496 -2 1872
rect 33 784 85 844
rect 549 424 601 484
rect 638 -604 692 -228
<< metal2 >>
rect -56 1872 -2 1882
rect -56 1378 -2 1496
rect -56 1371 2 1378
rect 635 1371 695 1380
rect -56 1369 92 1371
rect -56 1313 -54 1369
rect 2 1313 92 1369
rect -56 1311 92 1313
rect -56 1304 2 1311
rect -56 -32 -2 1304
rect 635 1302 695 1311
rect 33 844 85 854
rect 33 656 85 784
rect 33 604 601 656
rect 549 484 601 604
rect 549 414 601 424
rect -59 -41 1 -32
rect 638 -34 692 1302
rect -59 -110 1 -101
rect 635 -43 692 -34
rect 691 -99 692 -43
rect 635 -108 692 -99
rect 638 -228 692 -108
rect 638 -613 692 -604
<< via2 >>
rect -54 1313 2 1369
rect 635 1311 695 1371
rect -59 -101 1 -41
rect 635 -99 691 -43
<< metal3 >>
rect -59 1371 7 1374
rect 630 1371 700 1376
rect -59 1369 635 1371
rect -59 1313 -54 1369
rect 2 1313 635 1369
rect -59 1311 635 1313
rect 695 1311 700 1371
rect -59 1308 7 1311
rect 630 1306 700 1311
rect -64 -41 6 -36
rect 630 -41 696 -38
rect -64 -101 -59 -41
rect 1 -43 696 -41
rect 1 -99 635 -43
rect 691 -99 696 -43
rect 1 -101 696 -99
rect -64 -106 6 -101
rect 630 -104 696 -101
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729147637
transform 1 0 619 0 1 984
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729147637
transform 1 0 619 0 1 284
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729147637
transform 1 0 619 0 1 1684
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729147637
transform 1 0 619 0 1 -416
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729147637
transform 1 0 15 0 1 -416
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729147637
transform 1 0 15 0 1 284
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_9
timestamp 1729147637
transform 1 0 15 0 1 984
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_10
timestamp 1729147637
transform 1 0 15 0 1 1684
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729147637
transform 1 0 317 0 1 1684
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729147637
transform 1 0 317 0 1 984
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729147637
transform 1 0 317 0 1 284
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729147637
transform 1 0 317 0 1 -416
box -323 -300 323 300
<< labels >>
flabel metal3 1 -101 635 -41 0 FreeSans 320 0 0 0 D5
port 4 nsew
flabel metal2 549 484 601 656 0 FreeSans 160 0 0 0 D1
port 3 nsew
flabel poly 88 565 546 703 0 FreeSans 160 0 0 0 D2
port 6 nsew
flabel metal1 -58 -753 0 -697 0 FreeSans 480 0 0 0 VDD
port 8 nsew
<< end >>
